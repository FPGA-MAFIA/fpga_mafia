`include "macros.vh"

module d_mem_data_allignment
import big_core_pkg::*;
(
    


);



endmodule