modoule fifo_arb_TB();







endmodule

