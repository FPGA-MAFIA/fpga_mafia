package ps2_kbd_pkg;

parameter FIFO_WIDTH = 8;
parameter FIFO_DEPTH = 16;

endpackage