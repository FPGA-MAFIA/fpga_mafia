@00400000
A0 06 00 00 AC 06 00 00 B8 06 00 00 C4 06 00 00
D0 06 00 00 DC 06 00 00 E8 06 00 00 F4 06 00 00
00 07 00 00 0C 07 00 00 18 07 00 00 24 07 00 00
30 07 00 00 3C 07 00 00 48 07 00 00 48 45 4C 4C
4F 20 46 52 4F 4D 20 43 4F 52 45 20 31 20 54 48
52 45 41 44 20 50 4F 43 20 41 44 49 20 30 0A 00
20 20 20 20 00 00 00 00 48 45 4C 4C 4F 20 46 52
4F 4D 20 43 4F 52 45 20 31 20 54 48 52 45 41 44
20 31 0A 00 4D 41 54 52 49 58 20 31 0A 00 00 00
20 00 00 00 0A 00 00 00 0A 4D 41 54 52 49 58 20
32 0A 00 00 0A 4D 41 54 52 49 58 20 33 0A 00 00
01 00 00 00 02 00 00 00 03 00 00 00 04 00 00 00
05 00 00 00 06 00 00 00 07 00 00 00 08 00 00 00
09 00 00 00
@004000D4
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 3C 62 52 00 18 1C 1A 00 3C 42 40 00 3C 42 40
00 30 28 24 00 7E 02 3E 00 3C 42 02 00 7E 40 30
00 3C 42 42 00 3C 42 42 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 18 3C 66 00 1E 22 3E 00 3C 3E 02
00 1E 3E 22 00 7E 06 06 00 7E 06 06 00 3C 3E 02
00 66 66 66 00 7E 18 18 00 60 60 60 00 46 66 3E
00 06 06 06 00 42 66 5A 00 62 66 6E 00 3C 66 66
00 3E 66 66 00 3C 42 42 00 3E 66 66 00 7C 06 1E
00 7E 18 18 00 66 66 66 00 66 66 66 00 42 42 42
00 66 66 3C 00 66 66 3C 00 7E 20 10 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 18 18 1E 06 00 00 00 00 00 18 18 00
00 00 00 00 4A 46 3C 00 18 18 7E 00 3C 02 7E 00
38 42 3C 00 7E 20 20 00 40 42 3C 00 3E 42 3C 00
08 08 08 00 3C 42 3C 00 7C 40 3E 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 66 7E 66 00 3E 22 1E 00
02 3E 3C 00 22 3E 1E 00 7E 06 7E 00 7E 06 06 00
3A 22 3C 00 7E 66 66 00 18 18 7E 00 66 66 7C 00
3E 66 46 00 06 06 7E 00 5A 42 42 00 76 66 46 00
66 66 3C 00 3E 06 06 00 52 62 7C 00 3E 66 66 00
78 60 3E 00 18 18 18 00 66 7E 3C 00 66 3C 18 00
5A 7E 42 00 3C 66 66 00 18 18 18 00 08 04 7E 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 30 10 38 7C 30 10 38 38
30 10 38 38 30 10 38 7C 30 10 38 38 00 00 00 00
BA 48 84 82 78 AC 48 44 78 28 28 10 BA 38 10 28
7C 38 48 48 00 00 00 00
