delay(10);
random_gen_req(.trans(input_gen[NORTH]), .trans_valid(input_gen_valid[NORTH]) );
delay(1);
random_gen_req(.trans(input_gen[NORTH]), .trans_valid(input_gen_valid[NORTH]) );