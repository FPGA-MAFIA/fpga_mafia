@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 93 00 00 00 13 81 00 00 93 81 00 00
13 82 00 00 93 82 00 00 13 83 00 00 93 83 00 00
13 84 00 00 93 84 00 00 13 85 00 00 93 85 00 00
13 86 00 00 93 86 00 00 13 87 00 00 93 87 00 00
13 88 00 00 93 88 00 00 13 89 00 00 93 89 00 00
13 8A 00 00 93 8A 00 00 13 8B 00 00 93 8B 00 00
13 8C 00 00 93 8C 00 00 13 8D 00 00 93 8D 00 00
13 8E 00 00 93 8E 00 00 13 8F 00 00 93 8F 00 00
17 F1 01 00 13 01 01 F7 EF 00 80 0B 73 00 10 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
00 00 00 00 00 00 00 00 00 00 00 00 00 00 00 00
13 01 01 FE 23 2E 11 00 23 2C A1 00 23 2A B1 00
23 28 C1 00 23 26 D1 00 23 24 51 00 23 22 61 00
F3 22 90 00 93 82 12 00 73 90 92 00 83 20 C1 01
03 25 81 01 83 25 41 01 03 26 01 01 83 26 C1 00
83 22 81 00 03 23 41 00 13 01 01 02 73 00 20 30
13 01 01 FE 23 2E 81 00 13 04 01 02 93 07 10 00
23 26 F4 FE 83 27 C4 FE 93 87 17 00 23 26 F4 FE
6F F0 5F FF
