
`include "macros.vh"

module accel_core_mul_top 
import accel_core_pkg::*;
(
    input logic Clock,
    input logic Rst,
    
);
endmodule