ALIVE- NOT RELEVANT

