delay(1);  backdoor_fm_load();
//==========================================================
//  Randomly generate read/write requests
//==========================================================
// in this test will start with many write request to a small pull of addresses
// with a small delay between each request
// then will start with many read request to a small pull of addresses
// with a a big delay between each request - due to our missing stall functinality in the cache (after read miss)

create_addrs_pull(.local_num_tag_pull(10),//input
                  .local_num_set_pull(1),//input
                  .tag_pull(tag_pull),  //output
                  .set_pull(tag_pull)   //output
                  );

// send 50 wr request (Low Latency - B2B)
for(int i = 0; i<50; i++) begin
    random_wr(.local_min_req_delay(0), .local_max_req_delay(2));
end

// send 50 rd request (High Latency)
for(int i = 0; i<50; i++) begin
        random_rd(.local_min_req_delay(15), .local_max_req_delay(16));
end
