
//add here the alive tasks that you want to run