//First request
delay(10);
random_gen_req(.input_card(WEST));
//Second request
delay(10);
random_gen_req(.input_card(SOUTH)); 
delay(10);
random_gen_req(.input_card(SOUTH)); 