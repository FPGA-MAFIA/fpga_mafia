

fabric fabric (
.clk(clk),
.rst(rst)
);
