
`include "macros.vh"

module ifu_cache(


);
    

endmodule