package fabric_pkg;
`include "common_pkg.vh"

endpackage