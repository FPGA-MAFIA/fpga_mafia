parameter REQUESTS = 10;
