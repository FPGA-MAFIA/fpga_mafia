-	//
-	//File Name: fifo_arbiter.sv
-	//Description: The fifo_arbiter module.
-	//
-	module fifo_arbiter #(parameter int DATA_WIDTH=8,
-					parameter int FIFO_DEPTH=3,
-					parameter int NUM_CLIENTS=3)
-		(input			                  clk,
-		 input			                  rst,
-		 input [DATA_WIDTH-1:0]           din      [0:NUM_CLIENTS-1],
-		 input                            write    [NUM_CLIENTS-1:0],
-		 output                           full     [NUM_CLIENTS-1:0],
-		 output [$clog2(NUM_CLIENTS-1):0] src_num,           
-		 output                           valid,
-		 output [DATA_WIDTH-1:0]	      dout 
-		);
-	//INTERNAL VARIABLES
-	reg [DATA_WIDTH-1:0]     inside_din [0:NUM_CLIENTS-1];//maybe connect directly fifo to arbiter 
-	wire  [NUM_CLIENTS-1:0]	 ack;
-	logic                    empty [NUM_CLIENTS-1:0] ;
-	logic                    new_empty [NUM_CLIENTS-1:0];
-	
-	
-	
-	
-		arbiter #(.DATA_WIDTH(DATA_WIDTH),
-				.NUM_CLIENTS (NUM_CLIENTS))
-		arb
-			   (.clk(clk),
-			    .rst(rst),
-			    .req (new_empty),
-			    .din(inside_din),//get from fifo
-			    .src_num(src_num),
-			    .valid(valid),
-			    .ack(ack),
-			    .dout(dout)	);
-	genvar i;
-	generate
-		for (i=0; i<NUM_CLIENTS; i=i+1)begin
-			fifo #(.DATA_WIDTH(DATA_WIDTH),.FIFO_DEPTH(FIFO_DEPTH))
-				inside_fifo (.clk(clk),
-					     .rst(rst),
-					     .push(write[i]),
-					     .push_data(din[i]),
-					     .pop(ack[i]),
-					     .pop_data(inside_din[i]),
-					     .full(full[i]),
-					     .empty(empty[i]));//need to find how put !empty
-		end
-	endgenerate
-	
-	
-	
-	always @(posedge clk)
-	begin:NOT_EMPTY
-		for (int j=0; j<NUM_CLIENTS; j=j+1) begin
-			new_empty[j]=~empty[j];
-		end
-	end


endmodule: fifo_arbiter
