// this is the system verilog memory controller unit (MC)

module mc (
    input logic clk,
    input logic rst
)


//TODO create the memory controller unit

endmodule