module test ();
    initial $display("Hello, World!");
    initial $display("Hello again")
endmodule