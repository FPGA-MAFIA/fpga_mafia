//The fabric will instantiate a 3x3 mini_core_tile grid
