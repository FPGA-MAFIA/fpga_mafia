@00000000
13 00 00 00 13 00 00 00 13 00 00 00 13 00 00 00
13 00 00 00 6F 00 40 00 93 00 00 00 13 81 00 00
93 81 00 00 13 82 00 00 93 82 00 00 13 83 00 00
93 83 00 00 13 84 00 00 93 84 00 00 13 85 00 00
93 85 00 00 13 86 00 00 93 86 00 00 13 87 00 00
93 87 00 00 13 88 00 00 93 88 00 00 13 89 00 00
93 89 00 00 13 8A 00 00 93 8A 00 00 13 8B 00 00
93 8B 00 00 13 8C 00 00 93 8C 00 00 13 8D 00 00
93 8D 00 00 13 8E 00 00 93 8E 00 00 13 8F 00 00
93 8F 00 00 B7 02 C0 00 93 82 C2 00 03 A1 02 00
EF 00 90 5C 73 00 10 00
@000000A8
13 01 01 FD 23 26 81 02 13 04 01 03 93 07 05 00
23 2C B4 FC 23 2A C4 FC A3 0F F4 FC 03 27 84 FD
93 07 07 00 93 97 27 00 B3 87 E7 00 93 97 67 00
23 26 F4 FE 83 27 44 FD 93 97 27 00 23 24 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
B3 07 F7 00 23 22 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 93 87 07 14 B3 07 F7 00
23 20 F4 FE 83 47 F4 FD 37 07 40 00 13 07 47 0D
93 97 27 00 B3 07 F7 00 83 A7 07 00 13 87 07 00
83 27 44 FE 23 A0 E7 00 83 47 F4 FD 37 07 40 00
13 07 87 25 93 97 27 00 B3 07 F7 00 83 A7 07 00
13 87 07 00 83 27 04 FE 23 A0 E7 00 13 00 00 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 11 02 23 24 81 02 13 04 01 03 23 2E A4 FC
23 26 04 FE 23 24 04 FE 23 22 04 FE B7 07 C0 00
93 87 07 22 83 A7 07 00 23 22 F4 FE B7 07 C0 00
93 87 47 23 83 A7 07 00 23 24 F4 FE 6F 00 80 0B
83 27 C4 FE 03 27 C4 FD B3 07 F7 00 03 C7 07 00
93 07 A0 00 63 1A F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 6F 00 00 07 83 27 C4 FE 03 27 C4 FD
B3 07 F7 00 83 C7 07 00 03 27 84 FE 83 26 44 FE
13 86 06 00 93 05 07 00 13 85 07 00 EF F0 5F E8
83 27 44 FE 93 87 17 00 23 22 F4 FE 03 27 44 FE
93 07 00 05 63 12 F7 02 23 22 04 FE 83 27 84 FE
93 87 27 00 23 24 F4 FE 03 27 84 FE 93 07 80 07
63 14 F7 00 23 24 04 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 83 27 C4 FE 03 27 C4 FD B3 07 F7 00
83 C7 07 00 E3 9E 07 F2 B7 07 C0 00 93 87 07 22
03 27 44 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 84 FE 23 A0 E7 00 13 00 00 00 83 20 C1 02
03 24 81 02 13 01 01 03 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 2C B4 FC
23 2A C4 FC 03 27 84 FD 93 07 07 00 93 97 27 00
B3 87 E7 00 93 97 67 00 23 26 F4 FE 83 27 44 FD
93 97 27 00 23 24 F4 FE 03 27 84 FE 83 27 C4 FE
33 07 F7 00 B7 07 40 03 B3 07 F7 00 23 22 F4 FE
03 27 84 FE 83 27 C4 FE 33 07 F7 00 B7 07 40 03
93 87 07 14 B3 07 F7 00 23 20 F4 FE B7 07 40 00
13 87 C7 3D 83 27 C4 FD 93 97 27 00 B3 07 F7 00
83 A7 07 00 13 87 07 00 83 27 44 FE 23 A0 E7 00
B7 07 40 00 13 87 47 3F 83 27 C4 FD 93 97 27 00
B3 07 F7 00 83 A7 07 00 13 87 07 00 83 27 04 FE
23 A0 E7 00 13 00 00 00 03 24 C1 02 13 01 01 03
67 80 00 00 13 01 01 FE 23 2E 81 00 13 04 01 02
23 26 A4 FE 23 24 B4 FE B7 07 C0 00 93 87 07 22
03 27 84 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 C4 FE 23 A0 E7 00 13 00 00 00 03 24 C1 01
13 01 01 02 67 80 00 00 13 01 01 FE 23 2E 81 00
13 04 01 02 23 26 04 FE B7 07 40 03 23 24 F4 FE
23 26 04 FE 6F 00 40 02 83 27 C4 FE 93 97 27 00
03 27 84 FE B3 07 F7 00 23 A0 07 00 83 27 C4 FE
93 87 17 00 23 26 F4 FE 03 27 C4 FE B7 27 00 00
93 87 F7 57 E3 DA E7 FC 13 00 00 00 13 00 00 00
03 24 C1 01 13 01 01 02 67 80 00 00 13 01 01 FC
23 2E 11 02 23 2C 81 02 13 04 01 04 23 26 A4 FC
23 26 04 FE 23 24 04 FE 83 27 C4 FC 63 D6 07 02
83 27 C4 FE 13 87 17 00 23 26 E4 FE 13 07 04 FF
B3 07 F7 00 13 07 D0 02 23 80 E7 FE 83 27 C4 FC
B3 07 F0 40 23 26 F4 FC 83 27 C4 FC 93 05 A0 00
13 85 07 00 EF 00 D0 32 93 07 05 00 13 F7 F7 0F
83 27 C4 FE 93 86 17 00 23 26 D4 FE 13 07 07 03
13 77 F7 0F 93 06 04 FF B3 87 F6 00 23 80 E7 FE
83 27 C4 FC 93 05 A0 00 13 85 07 00 EF 00 10 27
93 07 05 00 23 26 F4 FC 83 27 C4 FC E3 46 F0 FA
23 24 04 FE 6F 00 00 07 83 27 84 FE 13 07 04 FF
B3 07 F7 00 83 C7 07 FE A3 0F F4 FC 03 27 C4 FE
83 27 84 FE B3 07 F7 40 93 87 F7 FF 13 07 04 FF
B3 07 F7 00 03 C7 07 FE 83 27 84 FE 93 06 04 FF
B3 87 F6 00 23 80 E7 FE 03 27 C4 FE 83 27 84 FE
B3 07 F7 40 93 87 F7 FF 13 07 04 FF B3 07 F7 00
03 47 F4 FD 23 80 E7 FE 83 27 84 FE 93 87 17 00
23 24 F4 FE 83 27 C4 FE 13 D7 F7 01 B3 07 F7 00
93 D7 17 40 13 87 07 00 83 27 84 FE E3 CE E7 F6
B7 07 C0 00 93 87 47 23 83 A7 07 00 23 22 F4 FE
B7 07 C0 00 93 87 07 22 83 A7 07 00 23 20 F4 FE
23 24 04 FE 6F 00 80 06 83 27 84 FE 13 07 04 FF
B3 07 F7 00 83 C7 07 FE 03 26 04 FE 83 25 44 FE
13 85 07 00 EF F0 DF B0 83 27 04 FE 93 87 17 00
23 20 F4 FE 03 27 04 FE 93 07 00 05 63 1A F7 00
23 20 04 FE 83 27 44 FE 93 87 27 00 23 22 F4 FE
03 27 44 FE 93 07 70 07 63 D4 E7 00 23 22 04 FE
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
83 27 C4 FE E3 4A F7 F8 B7 07 C0 00 93 87 07 22
03 27 04 FE 23 A0 E7 00 B7 07 C0 00 93 87 47 23
03 27 44 FE 23 A0 E7 00 13 00 00 00 83 20 C1 03
03 24 81 03 13 01 01 04 67 80 00 00 13 01 01 FD
23 26 81 02 13 04 01 03 23 2E A4 FC 23 26 04 FE
6F 00 00 01 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 83 27 C4 FD E3 46 F7 FE 13 00 00 00
13 00 00 00 03 24 C1 02 13 01 01 03 67 80 00 00
13 01 01 FD 23 26 81 02 13 04 01 03 23 2E A4 FC
03 27 C4 FD 93 07 E0 00 63 EA E7 0C 83 27 C4 FD
13 97 27 00 B7 07 40 00 93 87 07 00 B3 07 F7 00
83 A7 07 00 67 80 07 00 93 07 00 0C 23 26 F4 FE
6F 00 80 0B 93 07 90 0F 23 26 F4 FE 6F 00 C0 0A
93 07 40 0A 23 26 F4 FE 6F 00 00 0A 93 07 00 0B
23 26 F4 FE 6F 00 40 09 93 07 90 09 23 26 F4 FE
6F 00 80 08 93 07 20 09 23 26 F4 FE 6F 00 C0 07
93 07 20 08 23 26 F4 FE 6F 00 00 07 93 07 80 0F
23 26 F4 FE 6F 00 40 06 93 07 00 08 23 26 F4 FE
6F 00 80 05 93 07 00 09 23 26 F4 FE 6F 00 C0 04
93 07 80 08 23 26 F4 FE 6F 00 00 04 93 07 30 08
23 26 F4 FE 6F 00 40 03 93 07 60 0C 23 26 F4 FE
6F 00 80 02 93 07 10 0A 23 26 F4 FE 6F 00 C0 01
93 07 60 08 23 26 F4 FE 6F 00 00 01 93 07 00 08
23 26 F4 FE 13 00 00 00 83 27 C4 FE 13 85 07 00
03 24 C1 02 13 01 01 03 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 23 2A 91 00 13 04 01 02
23 26 A4 FE 83 27 C4 FE 93 05 A0 00 13 85 07 00
EF 00 10 01 93 07 05 00 B7 24 C0 03 13 85 07 00
EF F0 1F EC 93 07 05 00 23 A0 F4 00 83 27 C4 FE
93 05 A0 00 13 85 07 00 EF 00 40 76 93 07 05 00
93 05 A0 00 13 85 07 00 EF 00 80 7D 93 07 05 00
13 87 07 00 B7 27 C0 03 93 84 47 00 13 05 07 00
EF F0 1F E8 93 07 05 00 23 A0 F4 00 83 27 C4 FE
93 05 40 06 13 85 07 00 EF 00 40 72 93 07 05 00
93 05 A0 00 13 85 07 00 EF 00 80 79 93 07 05 00
13 87 07 00 B7 27 C0 03 93 84 87 00 13 05 07 00
EF F0 1F E4 93 07 05 00 23 A0 F4 00 83 27 C4 FE
93 05 80 3E 13 85 07 00 EF 00 40 6E 93 07 05 00
93 05 A0 00 13 85 07 00 EF 00 80 75 93 07 05 00
13 87 07 00 B7 27 C0 03 93 84 C7 00 13 05 07 00
EF F0 1F E0 93 07 05 00 23 A0 F4 00 03 27 C4 FE
B7 27 00 00 93 85 07 71 13 05 07 00 EF 00 00 6A
93 07 05 00 93 05 A0 00 13 85 07 00 EF 00 40 71
93 07 05 00 13 87 07 00 B7 27 C0 03 93 84 07 01
13 05 07 00 EF F0 DF DB 93 07 05 00 23 A0 F4 00
03 27 C4 FE B7 87 01 00 93 85 07 6A 13 05 07 00
EF 00 C0 65 93 07 05 00 93 05 A0 00 13 85 07 00
EF 00 00 6D 93 07 05 00 13 87 07 00 B7 27 C0 03
93 84 47 01 13 05 07 00 EF F0 9F D7 93 07 05 00
23 A0 F4 00 13 00 00 00 83 20 C1 01 03 24 81 01
83 24 41 01 13 01 01 02 67 80 00 00 13 01 01 FE
23 2E 11 00 23 2C 81 00 13 04 01 02 93 05 00 00
13 05 E0 01 EF F0 1F A5 B7 07 40 00 13 85 C7 03
EF F0 DF 83 23 26 04 FE 6F 00 C0 09 93 05 80 02
13 05 E0 01 EF F0 1F A3 03 25 C4 FE EF F0 1F AD
B7 27 C0 03 93 87 87 01 03 27 C4 FE 23 A0 E7 00
B7 27 C0 03 93 87 47 02 83 A7 07 00 23 22 F4 FE
93 05 20 03 13 05 E0 01 EF F0 DF 9F B7 07 40 00
13 85 07 06 EF F0 8F FE 93 05 20 03 13 05 E0 01
EF F0 5F 9E 03 25 44 FE EF F0 5F A8 03 25 C4 FE
EF F0 DF DC 23 24 04 FE 6F 00 00 01 83 27 84 FE
93 87 17 00 23 24 F4 FE 03 27 84 FE B7 27 00 00
93 87 F7 70 E3 D4 E7 FE 83 27 C4 FE 93 87 17 00
23 26 F4 FE 03 27 C4 FE B7 87 01 00 93 87 F7 69
E3 DE E7 F4 6F F0 9F F3 13 01 01 FF 23 26 11 00
23 24 81 00 13 04 01 01 93 05 00 00 13 05 80 02
EF F0 5F 97 B7 07 40 00 13 85 87 06 EF F0 0F F6
6F F0 9F FE 13 01 01 F6 23 2E 11 08 23 2C 81 08
23 2A 91 08 13 04 01 0A 93 05 00 00 13 05 60 04
EF F0 5F 94 B7 07 40 00 93 87 07 0B 03 A3 07 00
83 A8 47 00 03 A8 87 00 03 A5 C7 00 83 A5 07 01
03 A6 47 01 83 A6 87 01 03 A7 C7 01 83 A7 07 02
23 24 64 FA 23 26 14 FB 23 28 04 FB 23 2A A4 FA
23 2C B4 FA 23 2E C4 FA 23 20 D4 FC 23 22 E4 FC
23 24 F4 FC B7 07 40 00 93 87 07 0B 03 A3 07 00
83 A8 47 00 03 A8 87 00 03 A5 C7 00 83 A5 07 01
03 A6 47 01 83 A6 87 01 03 A7 C7 01 83 A7 07 02
23 22 64 F8 23 24 14 F9 23 26 04 F9 23 28 A4 F8
23 2A B4 F8 23 2C C4 F8 23 2E D4 F8 23 20 E4 FA
23 22 F4 FA 23 20 04 F6 23 22 04 F6 23 24 04 F6
23 26 04 F6 23 28 04 F6 23 2A 04 F6 23 2C 04 F6
23 2E 04 F6 23 20 04 F8 B7 07 40 00 13 85 47 08
EF F0 CF E6 23 26 04 FE 6F 00 80 07 23 24 04 FE
6F 00 C0 04 03 27 C4 FE 93 07 07 00 93 97 17 00
B3 87 E7 00 03 27 84 FE B3 87 E7 00 93 97 27 00
13 07 04 FF B3 07 F7 00 83 A7 87 FB 13 85 07 00
EF F0 DF 8D B7 07 40 00 13 85 07 09 EF F0 0F E2
83 27 84 FE 93 87 17 00 23 24 F4 FE 03 27 84 FE
93 07 20 00 E3 D8 E7 FA B7 07 40 00 13 85 47 09
EF F0 CF DF 83 27 C4 FE 93 87 17 00 23 26 F4 FE
03 27 C4 FE 93 07 20 00 E3 D2 E7 F8 B7 07 40 00
13 85 87 09 EF F0 8F DD 23 22 04 FE 6F 00 80 07
23 20 04 FE 6F 00 C0 04 03 27 44 FE 93 07 07 00
93 97 17 00 B3 87 E7 00 03 27 04 FE B3 87 E7 00
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 47 F9
13 85 07 00 EF F0 9F 84 B7 07 40 00 13 85 07 09
EF F0 CF D8 83 27 04 FE 93 87 17 00 23 20 F4 FE
03 27 04 FE 93 07 20 00 E3 D8 E7 FA B7 07 40 00
13 85 47 09 EF F0 8F D6 83 27 44 FE 93 87 17 00
23 22 F4 FE 03 27 44 FE 93 07 20 00 E3 D2 E7 F8
23 2E 04 FC 6F 00 40 10 23 2C 04 FC 6F 00 40 0E
23 2A 04 FC 6F 00 40 0C 03 27 C4 FD 93 07 07 00
93 97 17 00 B3 87 E7 00 03 27 84 FD B3 87 E7 00
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A4 07 F7
03 27 C4 FD 93 07 07 00 93 97 17 00 B3 87 E7 00
03 27 44 FD B3 87 E7 00 93 97 27 00 13 07 04 FF
B3 07 F7 00 83 A6 87 FB 03 27 44 FD 93 07 07 00
93 97 17 00 B3 87 E7 00 03 27 84 FD B3 87 E7 00
93 97 27 00 13 07 04 FF B3 07 F7 00 83 A7 47 F9
93 85 07 00 13 85 06 00 EF 00 00 24 93 07 05 00
B3 86 F4 00 03 27 C4 FD 93 07 07 00 93 97 17 00
B3 87 E7 00 03 27 84 FD B3 87 E7 00 93 97 27 00
13 07 04 FF B3 07 F7 00 23 A8 D7 F6 83 27 44 FD
93 87 17 00 23 2A F4 FC 03 27 44 FD 93 07 20 00
E3 DC E7 F2 83 27 84 FD 93 87 17 00 23 2C F4 FC
03 27 84 FD 93 07 20 00 E3 DC E7 F0 83 27 C4 FD
93 87 17 00 23 2E F4 FC 03 27 C4 FD 93 07 20 00
E3 DC E7 EE B7 07 40 00 13 85 47 0A EF F0 0F C3
23 28 04 FC 6F 00 80 07 23 26 04 FC 6F 00 C0 04
03 27 04 FD 93 07 07 00 93 97 17 00 B3 87 E7 00
03 27 C4 FC B3 87 E7 00 93 97 27 00 13 07 04 FF
B3 07 F7 00 83 A7 07 F7 13 85 07 00 EF F0 0F EA
B7 07 40 00 13 85 07 09 EF F0 4F BE 83 27 C4 FC
93 87 17 00 23 26 F4 FC 03 27 C4 FC 93 07 20 00
E3 D8 E7 FA B7 07 40 00 13 85 47 09 EF F0 0F BC
83 27 04 FD 93 87 17 00 23 28 F4 FC 03 27 04 FD
93 07 20 00 E3 D2 E7 F8 13 00 00 00 13 00 00 00
83 20 C1 09 03 24 81 09 83 24 41 09 13 01 01 0A
67 80 00 00 13 01 01 FD 23 26 11 02 23 24 81 02
13 04 01 03 23 2E A4 FC 23 26 04 FE 6F 00 00 05
83 27 C4 FD 93 97 27 00 93 05 80 02 13 85 07 00
EF F0 4F D6 03 25 C4 FE EF F0 4F E0 23 24 04 FE
6F 00 00 01 83 27 84 FE 93 87 17 00 23 24 F4 FE
03 27 84 FE B7 27 00 00 93 87 F7 70 E3 D4 E7 FE
83 27 C4 FE 93 87 17 00 23 26 F4 FE 03 27 C4 FE
B7 D7 9A 3B 93 87 F7 9F E3 D4 E7 FA 6F 00 00 00
13 01 01 FE 23 2E 11 00 23 2C 81 00 13 04 01 02
B7 07 C0 00 83 A7 07 00 23 26 F4 FE EF F0 CF D3
03 27 C4 FE 93 07 60 00 63 0E F7 02 03 27 C4 FE
93 07 60 00 63 CC E7 02 03 27 C4 FE 93 07 40 00
63 0A F7 00 03 27 C4 FE 93 07 50 00 63 08 F7 00
6F 00 C0 01 EF F0 9F A5 6F 00 80 01 EF F0 DF B2
6F 00 00 01 EF F0 1F B5 6F F0 DF FF 6F 00 00 00
03 27 C4 FE 93 07 40 00 63 04 F7 00 6F 00 00 00
93 07 00 00 13 85 07 00 83 20 C1 01 03 24 81 01
13 01 01 02 67 80 00 00 13 06 05 00 13 05 00 00
93 F6 15 00 63 84 06 00 33 05 C5 00 93 D5 15 00
13 16 16 00 E3 96 05 FE 67 80 00 00 63 40 05 06
63 C6 05 06 13 86 05 00 93 05 05 00 13 05 F0 FF
63 0C 06 02 93 06 10 00 63 7A B6 00 63 58 C0 00
13 16 16 00 93 96 16 00 E3 6A B6 FE 13 05 00 00
63 E6 C5 00 B3 85 C5 40 33 65 D5 00 93 D6 16 00
13 56 16 00 E3 96 06 FE 67 80 00 00 93 82 00 00
EF F0 5F FB 13 85 05 00 67 80 02 00 33 05 A0 40
63 48 B0 00 B3 05 B0 40 6F F0 DF F9 B3 05 B0 40
93 82 00 00 EF F0 1F F9 33 05 A0 40 67 80 02 00
93 82 00 00 63 CA 05 00 63 4C 05 00 EF F0 9F F7
13 85 05 00 67 80 02 00 B3 05 B0 40 E3 58 05 FE
33 05 A0 40 EF F0 1F F6 33 05 B0 40 67 80 02 00
