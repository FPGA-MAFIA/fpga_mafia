#1us;
$display("DONE COMPILATION AND ELABORATION");